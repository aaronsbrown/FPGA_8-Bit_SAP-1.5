module top (
    input clk,
    input rst_n,
    input usb_rx,
    output usb_tx,
    output [7:0] led
);
    
   

endmodule
