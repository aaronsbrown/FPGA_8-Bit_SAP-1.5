typedef struct packed {
    logic [3:0] opcode;
    logic [3:0] operand;
} instruction_t;

