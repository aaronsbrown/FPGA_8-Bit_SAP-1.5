module program_counter (
    input  wire clk,
    input  wire reset,
    // TODO: Add specific ports for program_counter
    input  wire [7:0] data_in,
    output wire [7:0] data_out
);

// TODO: Implement program_counter

endmodule
