module instruction_register (
    input  wire clk,
    input  wire reset,
    // TODO: Add specific ports for instruction_register
    input  wire [7:0] data_in,
    output wire [7:0] data_out
);

// TODO: Implement instruction_register

endmodule
