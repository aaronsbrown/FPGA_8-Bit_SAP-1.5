module alu (
    input  wire clk,
    input  wire reset,
    // TODO: Add specific ports for alu
    input  wire [7:0] data_in,
    output wire [7:0] data_out
);

// TODO: Implement alu

endmodule
