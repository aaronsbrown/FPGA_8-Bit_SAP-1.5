module ram (
    input  wire clk,
    input  wire reset,
    // TODO: Add specific ports for ram
    input  wire [7:0] data_in,
    output wire [7:0] data_out
);

// TODO: Implement ram

endmodule
