module eight_bit_fpga (
    // Define your module interface here
);
    // Your module implementation goes here
endmodule
